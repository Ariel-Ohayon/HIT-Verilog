//Behaviorial modeling Design.
//
//module Decoder3x8_ver1_Behave (D0,D1,D2,D3,D4,D5,D6,D7,A,B,C);
//output D0,D1,D2,D3,D4,D5,D6,D7;
//input  A,B,C;

